/* my_const.vh =  = = = = = = = = = = = = = = = = = = = = = = = = = = = *****
 **    basic constant definition					 ****
 ***       Ver. 1.0  2014.09.01						  ***
 ****									   **
 ***** (C) 2014 kimsyn (ET & VLSI system design labo. GCT ICE)  = = = = = = */


`define HIGH		1'b1
`define LOW  		1'b0

`define ON   		1'b1
`define OFF  		1'b0

`define YES  		1'b1
`define NO		1'b0

`define SET   		1'b1
`define RESET 		1'b0

`define ACTIVE  	1'b1
`define INACTIVE	1'b0

`define ACTIVE_N   	1'b0
`define INACTIVE_N 	1'b1

`define TRUE  	 	1'b1
`define FALSE 	 	1'b0

`define OK  		1'b1
`define NG  	 	1'b0

`define GOOD   	 	1'b1
`define NOGOOD 	 	1'b0

`define ERROR  	 	1'b1
`define NO_ERROR 	1'b0
