`default_nettype none

module ctrl_pla(
  input wire [3:0]    state,
  input wire [7:0]    instruction,
  input wire [2:0]    flag,
  output wire [17:0]  pla);

  assign pla = PLA(state, instruction, flag);

  //-- PLA function

  function [17:0] PLA;
    input [3:0] state;
    input [7:0] instruction;
    input [2:0] flag;
    begin
      casex({ state, instruction, flag})
        // instruction fetch
        15'b0000_XXXXXXXX_XXX : PLA = 18'b0_00_0_1_0100_01110_0000;
        15'b0001_XXXXXXXX_XXX : PLA = 18'b0_10_0_0_0000_00000_0100;
        15'b0010_XXXXXXXX_XXX : PLA = 18'b0_00_0_0_0111_00000_0101;
        //
        15'b0011_00000101_XXX : PLA = 18'b1_00_0_0_0001_00000_0001;
        15'b0011_00000110_XXX : PLA = 18'b1_00_0_0_0010_00000_0001;
        15'b0011_00000111_XXX : PLA = 18'b1_00_0_0_0011_00000_0001;
        15'b0011_00001001_XXX : PLA = 18'b1_00_0_0_0001_00000_0010;
        15'b0011_00001010_XXX : PLA = 18'b1_00_0_0_0010_00000_0010;
        15'b0011_00001011_XXX : PLA = 18'b1_00_0_0_0011_00000_0010;
        15'b0011_00001101_XXX : PLA = 18'b1_00_0_0_0001_00000_0011;
        15'b0011_00001110_XXX : PLA = 18'b1_00_0_0_0010_00000_0011;
        15'b0011_00001111_XXX : PLA = 18'b1_00_0_0_0011_00000_0011;
        15'b0011_100000XX_XXX : PLA = 18'b0_00_0_1_0100_01110_0000;
        15'b0100_100000XX_XXX : PLA = 18'b0_10_0_0_0000_00000_0100;
        15'b0101_100000XX_XXX : PLA = 18'b0_00_0_0_0100_00000_0101;
        15'b0110_100000XX_XXX : PLA = 18'b0_10_0_0_0000_00000_0000;
        15'b0111_10000001_XXX : PLA = 18'b1_00_0_0_0001_00000_0101;
        15'b0111_10000010_XXX : PLA = 18'b1_00_0_0_0010_00000_0101;
        15'b0111_10000011_XXX : PLA = 18'b1_00_0_0_0011_00000_0101;
        15'b0011_1010XX00_XXX : PLA = 18'b0_00_0_1_0100_01110_0000;
        15'b0100_1010XX00_XXX : PLA = 18'b0_10_0_0_0000_00000_0100;
        15'b0101_1010XX00_XXX : PLA = 18'b0_00_0_0_0100_00000_0101;
        15'b0110_10100100_XXX : PLA = 18'b0_00_0_0_0101_00000_0001;
        15'b0110_10101000_XXX : PLA = 18'b0_00_0_0_0101_00000_0010;
        15'b0110_10101100_XXX : PLA = 18'b0_00_0_0_0101_00000_0011;
        15'b0111_1010XX00_XXX : PLA = 18'b1_01_0_0_0000_00000_0000;
        15'b0011_001XXX01_XXX : PLA = 18'b0_00_0_0_0110_00000_0001;
        15'b0011_001XXX10_XXX : PLA = 18'b0_00_0_0_0110_00000_0010;
        15'b0011_001XXX11_XXX : PLA = 18'b0_00_0_0_0110_00000_0011;
        15'b0100_001000XX_XXX : PLA = 18'b0_00_1_1_0101_01000_0001;
        15'b0100_001001XX_XXX : PLA = 18'b0_00_1_1_0101_01010_0001;
        15'b0100_001010XX_XXX : PLA = 18'b0_00_1_1_0101_01011_0001;
        15'b0100_001011XX_XXX : PLA = 18'b0_00_1_1_0101_01101_0001;
        15'b0100_001100XX_XXX : PLA = 18'b0_00_1_1_0101_10000_0001;
        15'b0100_001101XX_XXX : PLA = 18'b0_00_1_1_0101_10001_0001;
        15'b0100_001111XX_XXX : PLA = 18'b0_00_1_1_0101_10010_0001;
        15'b0101_001XXXXX_XXX : PLA = 18'b1_00_0_0_0001_00000_0100;
        15'b0011_01000001_XXX : PLA = 18'b0_00_1_1_0110_01110_0001;
        15'b0011_01000010_XXX : PLA = 18'b0_00_1_1_0110_01110_0010;
        15'b0011_01000011_XXX : PLA = 18'b0_00_1_1_0110_01110_0011;
        15'b0011_01000101_XXX : PLA = 18'b0_00_1_1_0110_01111_0001;
        15'b0011_01000110_XXX : PLA = 18'b0_00_1_1_0110_01111_0010;
        15'b0011_01000111_XXX : PLA = 18'b0_00_1_1_0110_01111_0011;
        15'b0011_01010001_XXX : PLA = 18'b0_00_1_1_0110_10011_0001;
        15'b0011_01010010_XXX : PLA = 18'b0_00_1_1_0110_10011_0010;
        15'b0011_01010011_XXX : PLA = 18'b0_00_1_1_0110_10011_0011;
        15'b0100_010XXX01_XXX : PLA = 18'b1_00_0_0_0001_00000_0100;
        15'b0100_010XXX10_XXX : PLA = 18'b1_00_0_0_0010_00000_0100;
        15'b0100_010XXX11_XXX : PLA = 18'b1_00_0_0_0011_00000_0100;
        15'b0011_11000000_XXX : PLA = 18'b0_00_0_0_0100_00000_0000;
        15'b0100_11000000_XXX : PLA = 18'b0_10_0_0_0000_00000_0000;
        15'b0101_11000000_XXX : PLA = 18'b1_00_0_0_0000_00000_0101;
        15'b0011_11011XXX_XXX : PLA = 18'b0_00_0_1_0100_01110_0000;
        15'b0100_11011100_0XX : PLA = 18'b1_00_0_0_0000_00000_0100;
        15'b0100_11011100_1XX : PLA = 18'b0_10_0_0_0000_00000_0000;
        15'b0100_11011010_X0X : PLA = 18'b1_00_0_0_0000_00000_0100;
        15'b0100_11011010_X1X : PLA = 18'b0_10_0_0_0000_00000_0000;
        15'b0100_11011001_XX0 : PLA = 18'b1_00_0_0_0000_00000_0100;
        15'b0100_11011001_XX1 : PLA = 18'b0_10_0_0_0000_00000_0000;
        15'b0101_11011XXX_XXX : PLA = 18'b1_00_0_0_0000_00000_0101;
        15'b0011_00000000_XXX : PLA = 18'b0_00_0_0_0000_00000_0000;
        15'b0011_11111111_XXX : PLA = 18'b0_00_0_1_0000_01111_0000;
        15'b0100_11111111_XXX : PLA = 18'b1_00_0_0_0000_00000_0100;
        15'b0011_11101000_XXX : PLA = 18'b1_00_0_0_0000_00100_0000;
        15'b0011_11101001_XXX : PLA = 18'b1_00_0_0_0000_00101_0000;
        15'b0011_11101010_XXX : PLA = 18'b1_00_0_0_0000_00110_0000;
        //
        15'b0011_00000001_XXX : PLA = 18'b1_00_0_0_0001_00000_1000; // IN  ( IPORT -> A)
        15'b0011_00000100_XXX : PLA = 18'b1_00_0_0_1000_00000_0001; // OUT ( A -> OPORT)
        default : PLA = 18'bX_XX_X_X_XXXX_XXXXX_XXXX;
      endcase
    end
  endfunction

endmodule
